
module sigmoid
#(
    FLOAT_WIDTH = 31,
    LOG_FLOAT_WIDTH = 5
)
(
    input clk,
    input [FLOAT_WIDTH-1:0] x,

    output [FLOAT_WIDTH-1:0] y
);

    // ROM

    

    



endmodule
